library ieee;
use ieee.std_logic_1164.all;

entity invmixcolumn2 is 
    port (mi : in  std_logic_vector (31 downto 0);
          mo : out std_logic_vector (31 downto 0));
end entity;

architecture parallel of invmixcolumn2 is

    signal u      : std_logic_vector(31 downto 0);
    signal uu     : std_logic_vector(31 downto 0);
    signal uuu    : std_logic_vector(31 downto 0);
    signal uuuu   : std_logic_vector(31 downto 0);
    signal uuuuu  : std_logic_vector(31 downto 0);
    signal uuuuuu : std_logic_vector(31 downto 0);
    signal v      : std_logic_vector(31 downto 0);
    --signal y : std_logic_vector(31 downto 0);
    --signal t : std_logic_vector(59 downto 0);

begin
    
    proc : process(all)
      variable x, y : std_logic_vector(31 downto 0);
    begin
        
       x(7 downto 0)   := mi(31 downto 24);
       x(15 downto 8)  := mi(23 downto 16);
       x(23 downto 16) := mi(15 downto 8);
       x(31 downto 24) := mi(7  downto 0);

x(21) := x(21) xor x(5);
x(29) := x(29) xor x(21);
x(13) := x(13) xor x(29);
x(30) := x(30) xor x(14);
x(30) := x(30) xor x(13);
x(9) := x(9) xor x(17);
x(22) := x(22) xor x(13);
x(14) := x(14) xor x(22);
x(22) := x(22) xor x(6);
x(12) := x(12) xor x(20);
x(28) := x(28) xor x(12);
x(4) := x(4) xor x(28);
x(31) := x(31) xor x(23);
x(23) := x(23) xor x(30);
x(7) := x(7) xor x(23);
x(23) := x(23) xor x(15);
x(21) := x(21) xor x(4);
x(7) := x(7) xor x(22);
x(14) := x(14) xor x(21);
x(0) := x(0) xor x(23);
x(1) := x(1) xor x(9);
x(25) := x(25) xor x(1);
x(26) := x(26) xor x(10);
x(1) := x(1) xor x(0);
x(0) := x(0) xor x(24);
x(31) := x(31) xor x(22);
x(18) := x(18) xor x(2);
x(27) := x(27) xor x(7);
x(5) := x(5) xor x(13);
x(9) := x(9) xor x(8);
x(15) := x(15) xor x(14);
x(8) := x(8) xor x(23);
x(24) := x(24) xor x(7);
x(18) := x(18) xor x(25);
x(26) := x(26) xor x(25);
x(25) := x(25) xor x(9);
x(27) := x(27) xor x(18);
x(9) := x(9) xor x(24);
x(28) := x(28) xor x(23);
x(10) := x(10) xor x(9);
x(17) := x(17) xor x(16);
x(17) := x(17) xor x(31);
x(3) := x(3) xor x(11);
x(17) := x(17) xor x(25);    y(9) := x(17);
x(11) := x(11) xor x(26);
x(11) := x(11) xor x(27);
x(25) := x(25) xor x(1);    y(1) := x(25);
x(27) := x(27) xor x(19);
x(1) := x(1) xor x(24);    y(25) := x(1);
x(24) := x(24) xor x(16);
x(16) := x(16) xor x(0);    y(8) := x(16);
x(0) := x(0) xor x(8);
x(12) := x(12) xor x(11);
x(11) := x(11) xor x(23);
x(0) := x(0) xor x(31);    y(16) := x(0);
x(20) := x(20) xor x(31);
x(19) := x(19) xor x(11);
x(11) := x(11) xor x(31);
x(31) := x(31) xor x(15);    y(7) := x(31);
x(15) := x(15) xor x(7);    y(31) := x(15);
x(10) := x(10) xor x(18);    y(26) := x(10);
x(6) := x(6) xor x(14);
x(3) := x(3) xor x(18);
x(28) := x(28) xor x(3);    y(4) := x(28);
x(3) := x(3) xor x(7);
x(13) := x(13) xor x(21);
x(2) := x(2) xor x(25);
x(8) := x(8) xor x(24);    y(0) := x(8);
x(20) := x(20) xor x(27);
x(29) := x(29) xor x(12);    y(13) := x(29);
x(9) := x(9) xor x(17);    y(17) := x(9);
x(5) := x(5) xor x(20);
x(20) := x(20) xor x(4);    y(20) := x(20);
x(2) := x(2) xor x(17);
x(4) := x(4) xor x(12);
x(2) := x(2) xor x(26);    y(18) := x(2);
x(7) := x(7) xor x(31);    y(23) := x(7);
x(6) := x(6) xor x(29);
x(13) := x(13) xor x(29);    y(29) := x(13);
x(19) := x(19) xor x(10);
x(24) := x(24) xor x(0);    y(24) := x(24);
x(26) := x(26) xor x(10);    y(10) := x(26);
x(4) := x(4) xor x(28);    y(28) := x(4);
x(23) := x(23) xor x(7);    y(15) := x(23);
x(12) := x(12) xor x(20);    y(12) := x(12);
x(18) := x(18) xor x(2);    y(2) := x(18);
x(19) := x(19) xor x(2);    y(3) := x(19);
x(5) := x(5) xor x(4);    y(5) := x(5);
x(3) := x(3) xor x(19);    y(11) := x(3);
x(11) := x(11) xor x(3);    y(27) := x(11);
x(6) := x(6) xor x(5);    y(30) := x(6);
x(30) := x(30) xor x(6);    y(14) := x(30);
x(21) := x(21) xor x(5);    y(21) := x(21);
x(27) := x(27) xor x(11);    y(19) := x(27);
x(14) := x(14) xor x(30);    y(22) := x(14);
x(22) := x(22) xor x(14);    y(6) := x(22);


       --x(13) := x(13) xor x(29);
       --x(30) := x(30) xor x(14);
       --x(5) := x(5) xor x(13);
       --x(29) := x(29) xor x(21);
       --x(21) := x(21) xor x(5);
       --x(30) := x(30) xor x(21);
       --x(16) := x(16) xor x(0);
       --x(26) := x(26) xor x(10);
       --x(31) := x(31) xor x(30);
       --x(27) := x(27) xor x(3);
       --x(2) := x(2) xor x(26);
       --x(4) := x(4) xor x(20);
       --x(10) := x(10) xor x(18);
       --x(3) := x(3) xor x(19);
       --x(9) := x(9) xor x(17);
       --x(17) := x(17) xor x(25);
       --x(14) := x(14) xor x(6);
       --x(23) := x(23) xor x(30);
       --x(17) := x(17) xor x(16);
       --x(12) := x(12) xor x(4);
       --x(9) := x(9) xor x(1);
       --x(20) := x(20) xor x(28);
       --x(6) := x(6) xor x(22);
       --x(1) := x(1) xor x(0);
       --x(0) := x(0) xor x(24);
       --x(24) := x(24) xor x(16);
       --x(16) := x(16) xor x(8);
       --x(23) := x(23) xor x(15);
       --x(15) := x(15) xor x(31);
       --x(31) := x(31) xor x(7);
       --x(19) := x(19) xor x(27);
       --x(3) := x(3) xor x(2);
       --x(4) := x(4) xor x(31);
       --x(6) := x(6) xor x(21);
       --x(15) := x(15) xor x(6);
       --x(19) := x(19) xor x(23);
       --x(25) := x(25) xor x(9);
       --x(28) := x(28) xor x(12);
       --x(0) := x(0) xor x(15);
       --x(7) := x(7) xor x(15);
       --x(3) := x(3) xor x(18);
       --x(20) := x(20) xor x(3);
       --x(16) := x(16) xor x(31);    y(24) := x(16);
       --x(17) := x(17) xor x(15);
       --x(3) := x(3) xor x(31);
       --x(4) := x(4) xor x(11);
       --x(9) := x(9) xor x(31);
       --x(8) := x(8) xor x(23);
       --x(27) := x(27) xor x(15);
       --x(24) := x(24) xor x(23);    y(8) := x(24);
       --x(11) := x(11) xor x(3);
       --x(3) := x(3) xor x(23);
       --x(22) := x(22) xor x(30);
       --x(20) := x(20) xor x(15);
       --x(12) := x(12) xor x(31);
       --x(1) := x(1) xor x(8);
       --x(26) := x(26) xor x(25);
       --x(25) := x(25) xor x(1);    y(1) := x(25);
       --x(9) := x(9) xor x(0);    y(25) := x(9);
       --x(13) := x(13) xor x(28);
       --x(10) := x(10) xor x(1);
       --x(1) := x(1) xor x(17);    y(9) := x(1);
       --x(8) := x(8) xor x(0);    y(16) := x(8);
       --x(18) := x(18) xor x(26);
       --x(18) := x(18) xor x(17);    y(2) := x(18);
       --x(2) := x(2) xor x(17);    y(18) := x(2);
       --x(17) := x(17) xor x(9);    y(17) := x(17);
       --x(4) := x(4) xor x(19);
       --x(21) := x(21) xor x(13);
       --x(10) := x(10) xor x(17);
       --x(11) := x(11) xor x(10);    y(27) := x(11);
       --x(14) := x(14) xor x(21);
       --x(7) := x(7) xor x(14);    y(23) := x(7);
       --x(23) := x(23) xor x(7);    y(15) := x(23);
       --x(27) := x(27) xor x(26);
       --x(19) := x(19) xor x(10);    y(11) := x(19);
       --x(12) := x(12) xor x(27);    y(28) := x(12);
       --x(10) := x(10) xor x(2);    y(10) := x(10);
       --x(28) := x(28) xor x(4);
       --x(27) := x(27) xor x(11);    y(3) := x(27);
       --x(0) := x(0) xor x(16);    y(0) := x(0);
       --x(5) := x(5) xor x(20);    y(21) := x(5);
       --x(29) := x(29) xor x(4);
       --x(21) := x(21) xor x(5);    y(5) := x(21);
       --x(22) := x(22) xor x(29);    y(6) := x(22);
       --x(15) := x(15) xor x(23);    y(31) := x(15);
       --x(29) := x(29) xor x(5);    y(29) := x(29);
       --x(14) := x(14) xor x(22);    y(14) := x(14);
       --x(31) := x(31) xor x(15);    y(7) := x(31);
       --x(6) := x(6) xor x(22);    y(22) := x(6);
       --x(28) := x(28) xor x(12);    y(12) := x(28);
       --x(20) := x(20) xor x(12);    y(20) := x(20);
       --x(13) := x(13) xor x(29);    y(13) := x(13);
       --x(3) := x(3) xor x(27);    y(19) := x(3);
       --x(4) := x(4) xor x(20);    y(4) := x(4);
       --x(26) := x(26) xor x(10);    y(26) := x(26);
       --x(30) := x(30) xor x(14);    y(30) := x(30);

       mo(7 downto 0)   <= y(31 downto 24);
       mo(15 downto 8)  <= y(23 downto 16);
       mo(23 downto 16) <= y(15 downto 8);
       mo(31 downto 24) <= y(7  downto 0);

    end process;

end architecture;


